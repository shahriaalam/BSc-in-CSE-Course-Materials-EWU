* C:\Users\bmsha\OneDrive\Desktop\Project\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Mon May 22 00:45:02 2023



** Analysis setup **
.tran 0ns 5ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
